library verilog;
use verilog.vl_types.all;
entity MAGIC_BOX_vlg_vec_tst is
end MAGIC_BOX_vlg_vec_tst;
