library verilog;
use verilog.vl_types.all;
entity Magic_Box_vlg_vec_tst is
end Magic_Box_vlg_vec_tst;
