library verilog;
use verilog.vl_types.all;
entity COUNTER_LPM_vlg_vec_tst is
end COUNTER_LPM_vlg_vec_tst;
