library verilog;
use verilog.vl_types.all;
entity all_uart_vlg_vec_tst is
end all_uart_vlg_vec_tst;
